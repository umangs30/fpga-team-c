module storage();
reg [7:0] a[8:0][0:2];
assign a[0][0]=0;
assign a[0][1]=0;
assign 
assign a[1][0]=1;
assign a[1][1]=0;
//16
assign a[2][0]=1;
assign a[2][1]=2;
//91
assign a[3][0]=1;
assign a[3][1]=2;
//
assign a[4][0]=4;
assign a[4][1]=0;
//58
assign a[5][0]=4;
assign a[5][1]=2;

assign a[6][0]=5;
assign a[6][1]=6;

assign a[7][0]=6;
assign a[7][1]=6;

assign a[8][0]=7;
assign a[8][1]=8;



